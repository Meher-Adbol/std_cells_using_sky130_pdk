VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO and2b
  CLASS BLOCK ;
  FOREIGN and2b ;
  ORIGIN 1.750 0.350 ;
  SIZE 10.230 BY 3.020 ;
  OBS
      LAYER nwell ;
        RECT -1.470 0.720 0.380 2.350 ;
        RECT 1.670 0.920 3.880 2.550 ;
        RECT 6.630 0.720 8.480 2.350 ;
        RECT -1.470 0.710 -0.250 0.720 ;
        RECT 6.630 0.710 7.850 0.720 ;
      LAYER li1 ;
        RECT -1.290 2.170 -0.940 2.670 ;
        RECT 1.850 2.370 2.150 2.670 ;
        RECT -1.290 0.900 -0.270 2.170 ;
        RECT -0.080 0.900 0.200 2.170 ;
        RECT 1.850 1.100 2.780 2.370 ;
        RECT 2.970 1.100 3.230 2.370 ;
        RECT 3.420 1.100 3.700 2.670 ;
        RECT 6.810 2.170 7.160 2.670 ;
        RECT 3.950 1.300 4.850 1.700 ;
        RECT 4.600 0.920 4.940 1.100 ;
        RECT 0.000 0.720 0.200 0.900 ;
        RECT 0.650 0.720 1.000 0.820 ;
        RECT 1.430 0.750 4.940 0.920 ;
        RECT 6.810 0.900 7.830 2.170 ;
        RECT 8.020 0.900 8.300 2.170 ;
        RECT 1.430 0.720 1.610 0.750 ;
        RECT 0.000 0.550 1.610 0.720 ;
        RECT 8.100 0.720 8.300 0.900 ;
        RECT 0.000 0.370 0.200 0.550 ;
        RECT 0.650 0.450 1.000 0.550 ;
        RECT -0.950 -0.050 -0.270 0.370 ;
        RECT -0.080 -0.050 0.200 0.370 ;
        RECT 2.100 0.150 2.780 0.570 ;
        RECT 2.970 0.150 3.230 0.570 ;
        RECT 3.420 0.150 4.680 0.570 ;
        RECT 4.870 0.150 5.130 0.570 ;
        RECT 5.320 0.150 6.000 0.570 ;
        RECT 8.100 0.550 8.480 0.720 ;
        RECT 8.100 0.370 8.300 0.550 ;
        RECT -0.950 -0.350 -0.550 -0.050 ;
        RECT 2.100 -0.350 2.500 0.150 ;
        RECT 3.000 -0.150 3.200 0.150 ;
        RECT 4.900 -0.150 5.100 0.150 ;
        RECT 3.000 -0.350 5.100 -0.150 ;
        RECT 5.600 -0.350 6.000 0.150 ;
        RECT 7.150 -0.050 7.830 0.370 ;
        RECT 8.020 -0.050 8.300 0.370 ;
        RECT 7.150 -0.350 7.550 -0.050 ;
      LAYER met1 ;
        RECT -1.750 2.370 8.480 2.670 ;
        RECT 3.950 1.450 4.250 1.700 ;
        RECT 2.950 1.300 4.250 1.450 ;
        RECT 2.950 1.150 4.200 1.300 ;
        RECT 3.850 0.150 4.200 1.150 ;
        RECT -1.750 -0.350 8.480 -0.050 ;
  END
END and2b
END LIBRARY

