VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 3_input_NAND_wload
  CLASS BLOCK ;
  FOREIGN 3_input_NAND_wload ;
  ORIGIN 7.480 -0.270 ;
  SIZE 11.130 BY 3.030 ;
  PIN Ain
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT -7.480 1.420 -7.030 1.720 ;
    END
  END Ain
  PIN Abar
    ANTENNAGATEAREA 0.378000 ;
    ANTENNADIFFAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT -5.950 1.520 -5.710 2.860 ;
        RECT -5.950 1.350 -5.190 1.520 ;
        RECT -5.950 1.180 -5.710 1.350 ;
        RECT -5.360 1.340 -5.190 1.350 ;
        RECT -5.970 0.810 -5.690 1.180 ;
        RECT -5.360 0.980 -5.000 1.340 ;
    END
  END Abar
  PIN Bin
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT -5.520 2.140 -5.160 2.500 ;
    END
  END Bin
  PIN Cin
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 0.930 1.230 1.290 1.590 ;
    END
  END Cin
  PIN Y
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 1.176000 ;
    PORT
      LAYER li1 ;
        RECT -2.530 2.660 -0.160 2.830 ;
        RECT -2.530 2.420 -2.360 2.660 ;
        RECT -1.440 2.420 -1.260 2.660 ;
        RECT -0.340 2.420 -0.160 2.660 ;
        RECT -4.830 2.030 -4.460 2.420 ;
        RECT -3.730 2.030 -3.370 2.420 ;
        RECT -2.630 2.030 -2.270 2.420 ;
        RECT -1.530 2.030 -1.170 2.420 ;
        RECT -0.430 2.030 -0.070 2.420 ;
        RECT -4.740 1.410 -4.560 2.030 ;
        RECT -3.640 1.410 -3.460 2.030 ;
        RECT -1.440 1.410 -1.260 2.030 ;
        RECT 1.500 1.420 1.840 1.720 ;
        RECT -4.740 1.240 -1.260 1.410 ;
        RECT -4.740 1.000 -4.560 1.240 ;
        RECT -3.640 1.000 -3.460 1.240 ;
        RECT -1.460 1.180 -1.260 1.240 ;
        RECT -4.830 0.700 -4.470 1.000 ;
        RECT -3.730 0.700 -3.370 1.000 ;
      LAYER met1 ;
        RECT 1.500 1.400 1.840 1.720 ;
        RECT -1.500 1.160 1.840 1.400 ;
    END
  END Y
  PIN Ybar
    ANTENNADIFFAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 2.920 1.520 3.160 2.860 ;
        RECT 2.920 1.350 3.620 1.520 ;
        RECT 2.920 1.180 3.160 1.350 ;
        RECT 2.900 0.810 3.180 1.180 ;
    END
  END Ybar
  OBS
      LAYER nwell ;
        RECT -6.970 2.660 -5.500 3.160 ;
        RECT 1.900 2.660 3.370 3.160 ;
        RECT -6.970 1.820 3.370 2.660 ;
        RECT -6.970 1.540 -5.500 1.820 ;
        RECT 1.900 1.540 3.370 1.820 ;
      LAYER li1 ;
        RECT -6.910 3.230 3.370 3.240 ;
        RECT -6.950 3.040 3.370 3.230 ;
        RECT -6.950 3.030 -6.720 3.040 ;
        RECT -6.550 3.030 3.370 3.040 ;
        RECT -6.370 2.860 -6.200 3.030 ;
        RECT -6.800 1.800 -6.160 2.860 ;
        RECT -4.190 2.420 -4.010 3.030 ;
        RECT -3.090 2.440 -2.910 3.030 ;
        RECT -4.280 2.030 -3.920 2.420 ;
        RECT -3.180 2.030 -2.820 2.440 ;
        RECT 0.210 2.420 0.390 3.030 ;
        RECT 2.500 2.860 2.670 3.030 ;
        RECT -2.080 2.030 -1.720 2.420 ;
        RECT -0.980 2.030 -0.620 2.420 ;
        RECT 0.120 2.030 0.900 2.420 ;
        RECT -3.090 1.760 -2.910 2.030 ;
        RECT -1.990 1.760 -1.810 2.030 ;
        RECT -3.090 1.580 -1.810 1.760 ;
        RECT -0.890 1.760 -0.710 2.030 ;
        RECT 0.200 1.760 0.400 2.030 ;
        RECT 2.070 1.800 2.710 2.860 ;
        RECT -0.890 1.580 0.400 1.760 ;
        RECT -6.810 0.810 -6.140 1.180 ;
        RECT -6.360 0.520 -6.190 0.810 ;
        RECT -4.280 0.700 -3.920 1.000 ;
        RECT -3.180 0.700 -2.820 1.000 ;
        RECT -2.630 0.700 -2.270 1.000 ;
        RECT -2.070 0.700 -1.710 1.000 ;
        RECT -1.520 0.700 -1.160 1.000 ;
        RECT -0.970 0.700 -0.610 1.000 ;
        RECT -0.430 0.700 -0.070 1.000 ;
        RECT 0.120 0.700 0.890 1.000 ;
        RECT 2.060 0.810 2.730 1.180 ;
        RECT -0.880 0.520 -0.700 0.700 ;
        RECT 0.210 0.690 0.890 0.700 ;
        RECT 0.210 0.520 0.390 0.690 ;
        RECT 2.510 0.520 2.680 0.810 ;
        RECT -6.940 0.320 3.650 0.520 ;
      LAYER met1 ;
        RECT -6.950 2.980 3.650 3.300 ;
        RECT -3.110 1.760 -2.890 2.980 ;
        RECT -2.040 1.760 -1.750 1.790 ;
        RECT -3.110 1.580 -1.750 1.760 ;
        RECT -2.040 1.550 -1.750 1.580 ;
        RECT -0.950 1.760 -0.660 1.790 ;
        RECT 0.180 1.760 0.420 2.980 ;
        RECT -0.950 1.580 0.420 1.760 ;
        RECT -0.950 1.550 -0.660 1.580 ;
        RECT -6.950 0.270 3.650 0.570 ;
  END
END 3_input_NAND_wload
END LIBRARY

