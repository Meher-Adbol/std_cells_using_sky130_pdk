* EE671 VLSI Design - Course Project 01 Group 12
* Name: Aditya Tare (24M1169), Gautam Govindaraju (24M1166), Ritoo Verma (24M1185), Sachin Soneria (24M1178)
* D flip flop (Negative Edge triggered)

*Including sky130 device model
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* Power supply
Vdd vdd gnd DC 1.8

* Input signals
* Vdin din gnd pulse(0 1.8 2.5ns 60ps 60ps 10ns 20ns)
* Vclk clock gnd pulse(0 1.8 0 10ps 10ps 5ns 10ns)
* Vdin din gnd pulse(0 1.8 4774ps 60ps 60ps 10ns 20ns) 	; Setup Time
* Vclk clock gnd pulse(0 1.8 0 10ps 10ps 5ns 10ns)	; Setup Time
* Vdin din gnd pulse(0 1.8 5.92ns 10ps 10ps 8ns 16ns) 	; Hold Time
* Vclk clock gnd pulse(0 1.8 5ns 10ps 10ps 5ns 10ns)  	; Hold Time
Vdin din gnd pulse(0 1.8 4198ps 1000ps 1000ps 8ns 16ns) 	; Library File
Vclk clock gnd pulse(0 1.8 0ps 10ps 10ps 5ns 10ns)  	; Library File

* Defining Subcircuit of Negative Edge Triggered DFF
.subckt dff D clk Q vdd gnd

X0 Dbar D vdd vdd sky130_fd_pr__pfet_01v8 ad=0.441 pd=3.22 as=0.378 ps=3.12 w=1.26 l=0.15
X1 Dbar D gnd gnd sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.126 ps=1.44 w=0.42 l=0.15
X2 2 1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.441 pd=3.22 as=0.378 ps=3.12 w=1.26 l=0.15
X3 2 1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.126 ps=1.44 w=0.42 l=0.15
X4 clk_inv clk vdd vdd sky130_fd_pr__pfet_01v8 ad=0.378 pd=3.12 as=0.378 ps=3.12 w=1.26 l=0.15
X5 clk_inv clk gnd gnd sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X6 3 2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.441 pd=3.22 as=0.378 ps=3.12 w=1.26 l=0.15
X7 3 2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.126 ps=1.44 w=0.42 l=0.15
X8 Qin 4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.378 pd=3.12 as=0.378 ps=3.12 w=1.26 l=0.15
X9 Qin 4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X10 5 Qin vdd vdd sky130_fd_pr__pfet_01v8 ad=0.441 pd=3.22 as=0.378 ps=3.12 w=1.26 l=0.15
X11 5 Qin gnd gnd sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.126 ps=1.44 w=0.42 l=0.15
X12 Q Qin vdd vdd sky130_fd_pr__pfet_01v8 ad=0.378 pd=3.12 as=0.378 ps=3.12 w=1.26 l=0.15
X13 Q Qin gnd gnd sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X14 3 clk 1 vdd sky130_fd_pr__pfet_01v8 ad=0.441 pd=3.22 as=0.504 ps=3.32 w=1.26 l=0.15
X15 3 clk_inv 1 gnd sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X16 5 clk_inv 4 vdd sky130_fd_pr__pfet_01v8 ad=0.441 pd=3.22 as=0.504 ps=3.32 w=1.26 l=0.15
X17 5 clk 4 gnd sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X18 2 clk 4 vdd sky130_fd_pr__pfet_01v8 ad=0.441 pd=3.22 as=0.504 ps=3.32 w=1.26 l=0.15
X19 2 clk_inv 4 gnd sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15
X20 Dbar clk_inv 1 vdd sky130_fd_pr__pfet_01v8 ad=0.441 pd=3.22 as=0.504 ps=3.32 w=1.26 l=0.15
X21 Dbar clk 1 gnd sky130_fd_pr__nfet_01v8 ad=0.147 pd=1.54 as=0.168 ps=1.64 w=0.42 l=0.15

C0 1 clk 0.076351f
C1 4 Q 0.002729f
C2 4 Qin 0.182473f
C3 4 clk_inv 0.867807f
C4 gnd D 1.35e-19
C5 clk Dbar 0.069862f
C6 clk 3 0.081248f
C7 2 5 2.86e-20
C8 2 clk 0.123158f
C9 1 Qin 2.33e-20
C10 1 clk_inv 0.976341f
C11 clk 5 0.013526f
C12 4 vdd 0.530653f
C13 Dbar clk_inv 0.279964f
C14 Qin 3 2.7e-20
C15 clk_inv 3 0.180625f
C16 1 D 6.61e-20
C17 2 Qin 0.002024f
C18 2 clk_inv 0.402873f
C19 Dbar D 0.038014f
C20 1 vdd 0.514643f
C21 5 Qin 0.169497f
C22 clk_inv 5 0.151278f
C23 Q clk 3.69e-20
C24 2 D 9.02e-21
C25 clk Qin 0.039507f
C26 clk clk_inv 0.24915f
C27 Dbar vdd 0.438696f
C28 4 gnd 1.158879f
C29 vdd 3 0.232927f
C30 2 vdd 1.213519f
C31 clk D 0.008498f
C32 vdd 5 0.262206f
C33 Q Qin 0.035751f
C34 Q clk_inv 2.49e-19
C35 clk vdd 1.14327f
C36 clk_inv Qin 0.258663f
C37 1 gnd 1.012704f
C38 4 1 0.004918f
C39 gnd Dbar 0.170931f
C40 gnd 3 0.037234f
C41 D clk_inv 1.67e-19
C42 2 gnd 0.059469f
C43 4 3 1.1e-20
C44 Q vdd 0.132627f
C45 vdd Qin 1.128015f
C46 vdd clk_inv 1.298286f
C47 2 4 0.152494f
C48 gnd 5 0.039708f
C49 gnd clk 0.34179f
C50 4 5 0.19776f
C51 D vdd 0.122108f
C52 4 clk 0.112107f
C53 1 Dbar 0.156332f
C54 1 3 0.187673f
C55 2 1 0.127121f
C56 Dbar 3 3.19e-19
C57 2 Dbar 0.003951f
C58 gnd Qin 0.056289f
C59 gnd clk_inv 0.469403f
C60 2 3 0.155633f
C61 gnd 0 1.130442f
C62 clk 0 2.35632f
C63 4 0 0.361989f
C64 1 0 0.322242f
C65 vdd 0 7.203994f
C66 Q 0 0.156718f
C67 5 0 0.115382f
C68 Qin 0 0.556712f
C69 3 0 0.101442f
C70 clk_inv 0 1.028028f
C71 2 0 0.344999f
C72 Dbar 0 0.152824f
C73 D 0 0.316317f
.ends dff

* Instantiating Subcircuit of D Flip flop
Xdff1 din clock out vdd gnd dff

* Transient Analysis
.tran 0.1ns 50ns 0 100ps

.control
run

meas tran tr TRIG v(out) VAL = 0.36 RISE = 1 TARG v(out) VAL = 1.44 RISE = 1
meas tran tf TRIG v(out) VAL = 1.44 FALL = 1 TARG v(out) VAL = 0.36 FALL = 2
meas tran tplh TRIG v(clock) VAL = 0.9 FALL = 1 TARG v(out) VAL = 0.9 RISE = 2
meas tran tphl TRIG v(clock) VAL = 0.9 FALL = 2 TARG v(out) VAL = 0.9 FALL = 2

let delta = abs(tr - tf)

let tprop = (tplh + tphl)/2

*meas tran tset TRIG v(din) VAL = 0.9 FALL = 1 TARG v(clock) VAL = 0.9 FALL = 2
*meas tran tset TRIG v(din) VAL = 0.9 RISE = 1 TARG v(clock) VAL = 0.9 FALL = 1
meas tran thold TRIG v(clock) VAL = 0.9 FALL = 1 TARG v(din) VAL = 0.9 RISE = 1

print tr
print tf
print delta
print tprop
*print tset
print thold

set color0=white
set color1=black
set color2=blue
set color3=purple
set color4=red
set xbrushwidth=5

plot out din+3  clock+6

.endc
.end