
* SkyWater PDK
* simple inverter

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* Voltage Sources:

Vdd vdd gnd DC 1.8
V1 in gnd PULSE(0 1.8 0 1000p 1000p 1n 6n)

* Subcircuit of inverter

.subckt not1 a vdd vss z
X0 z a vss vss sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.126 ps=1.44 w=0.42 l=0.15
X1 z a vdd vdd sky130_fd_pr__pfet_01v8 ad=0.378 pd=3.12 as=0.378 ps=3.12 w=1.26 l=0.15 

** Capacitors from PEX **

* C0 z vdd 0.130174f
* C1 a z 0.033116f
* C2 a vdd 0.108028f
* C3 z vss 0.171025f
* C4 a vss 0.33541f
* C5 vdd vss 0.529498f

.ends

* Instantiating Inverter with Load Capacitor or Inverter
Xnot1 in vdd gnd out not1
*Xnot2 out vdd gnd out2 not1

* Cload out gnd 100f


*Simulation Command:

.tran 1ps 10ns 0 10p
.control


******************** CONTROL STRUCTURE ********************

set color0=white
set color1=black
set color2=red
set color3=blue
set color4=green
run
meas tran Ipeak_rise MAX I(Vdd) from=0 to=1000p
meas tran Ipeak_fall MIN I(Vdd) from=2000e-12 to=3000e-12
let RISE_POWER= (0.5 * 10e-12 * Ipeak_rise *1.8)/3000e-12
let FALL_POWER= (0.5 * 10e-12 * Ipeak_fall * 1.8)/3000e-12
print RISE_POWER
print FALL_POWER
set xbrushwidth=4
plot I(V1) V(in)

******************** STATIC POWER CHARACTERISTICS ********************

* let StaticPower = I(Vdd) * Vdd
* print StaticPower

******************** DYNAMIC POWER CHARACTERISTICS ********************
* In this For loop we are changing values of Cload and Input Slew through variables 'val' and 'varx' respectively.
* we are measuring the peak value of current on rising and falling edge of the input voltage , this value is used to measure dynamic power.

* foreach val 0.5e-15 10e-15 100e-15
	* foreach varx 10e-12 100e-12 1000e-12
		* let a1=0
		* let a2=$varx
		* let b1=(3000e-12 - $varx)
		* let b2=(3000e-12)
		* let hold=(3000e-12 - 2 * $varx)
        * alter @Cload $val
		* alter @V1[PULSE] [ 0 1.8 0 $varx $varx $&hold 6n ]
		* echo CLoad is $val InputSlew is $varx
		* echo rise from 0 to $&a2
		* echo fall from $&b1 to $&b2
		* run	
		* meas tran Ipeak_rise MAX I(Vdd) from=0 to=$&a2
		* meas tran Ipeak_fall MIN I(Vdd) from=$&b1 to=$&b2
		* let RISE_POWER= (0.5* $varx * Ipeak_rise *1.8)/$&b2
		* let FALL_POWER= (0.5 *$varx * Ipeak_fall * 1.8)/$&b2
		* print RISE_POWER
		* print FALL_POWER
		* reset
	* end	
* end



******************** TIMING CHARACTERISTICS ********************
* In this For loop we are changing values of Cload and Input Slew through variables 'val' and 'varx' respectively.
* we are measuring the time for rising and falling edges of the output

* foreach val 0.5e-15 10e-15 100e-15
	* foreach varx 10e-12 100e-12 1000e-12
        * alter @Cload $val
		* alter @V1[PULSE] [ 0 1.8 0 $varx $varx 3n 6n ]
		* echo CLoad is $val InputSlew is $varx
		* run
		* meas tran T_RISE TRIG v(out) VAL = 0.36 RISE = 1 TARG v(out) VAL = 1.44 RISE = 1
		* meas tran T_FALL TRIG v(out) VAL = 1.44 FALL = 1 TARG v(out) VAL = 0.36 FALL = 1
		* meas tran CELL_RISE_DELAY TRIG v(in)  VAL = 0.9 FALL = 1 TARG v(out) VAL = 0.9 RISE = 1
		* meas tran CELL_FALL_DELAY TRIG v(in)  VAL = 0.9 RISE = 1 TARG v(out) VAL = 0.9 FALL = 1		
		* reset
	* end	
* end




******************** INPUT CAPACITANCE ********************
* In this part we first inject a known voltage source and we integrate the current during falling and rising edges of the voltage source , these values
* of current are used to calculate input capacitance.
 

*meas tran I_integ_rise INTEG I(V1) from=0p to =500p
*meas tran I_integ_fall INTEG I(V1) from=1500p to =2000p
*let InputCapRise=I_integ_rise/1.8
*let InputCapFall=I_integ_fall/1.8
*let Avg_Cap=(InputCapRise+InputCapFall)/2
*print InputCapRise InputCapFall Avg_Cap



.endc
