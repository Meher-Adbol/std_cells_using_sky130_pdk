magic
tech sky130A
timestamp 1726337622
<< nwell >>
rect -510 244 1916 252
rect -510 232 1209 244
rect -510 229 -504 232
rect -486 231 -467 232
rect -363 229 -268 232
rect -249 231 -230 232
rect -127 231 173 232
rect 192 231 211 232
rect -363 102 -274 229
rect -369 82 -274 102
rect -127 222 -76 231
rect 95 229 173 231
rect -127 218 -18 222
rect -127 82 -76 218
rect 95 70 167 229
rect 313 82 353 232
rect 377 231 396 232
rect 490 231 1209 232
rect 490 229 1130 231
rect 1136 229 1209 231
rect 490 222 1123 229
rect 490 217 631 222
rect 490 215 632 217
rect 500 82 580 215
rect 744 76 808 222
rect 951 82 1123 222
rect 1136 82 1203 229
rect 1270 173 1310 244
rect 1320 236 1795 244
rect 1320 232 1348 236
rect 1457 232 1795 236
rect 1320 231 1353 232
rect 1457 231 1811 232
rect 1267 165 1312 173
rect 1320 165 1348 231
rect 1457 222 1575 231
rect 1601 222 1631 231
rect 1729 229 1795 231
rect 1457 165 1558 222
rect 1729 165 1787 229
rect 1267 133 1787 165
rect 1270 82 1310 133
rect 1320 82 1348 133
rect 1457 82 1558 133
rect 1729 82 1787 133
rect 767 70 886 76
rect 951 70 1009 82
rect 1747 70 1781 82
<< poly >>
rect -100 222 -3 237
rect 325 234 452 249
rect -100 74 -85 222
rect 327 181 342 234
rect 490 222 1017 237
rect 316 173 352 181
rect 316 153 324 173
rect 344 153 352 173
rect 316 145 352 153
rect -112 66 -76 74
rect -112 46 -104 66
rect -84 46 -76 66
rect -112 38 -76 46
rect -190 -28 -175 -7
rect -18 -28 -3 -18
rect 490 -28 505 222
rect 761 74 797 82
rect 533 66 569 74
rect 533 46 541 66
rect 561 46 569 66
rect 761 54 769 74
rect 789 54 797 74
rect 761 46 797 54
rect 533 38 569 46
rect -190 -43 505 -28
rect 554 -14 569 38
rect 763 -14 778 46
rect 554 -15 631 -14
rect 554 -29 646 -15
rect 763 -29 881 -14
rect 1002 -28 1017 222
rect 1485 222 1631 237
rect 1270 156 1304 163
rect 1270 138 1278 156
rect 1296 138 1304 156
rect 1270 133 1304 138
rect 1279 100 1294 133
rect 1485 74 1500 222
rect 1474 66 1510 74
rect 1747 70 1781 100
rect 1474 46 1482 66
rect 1502 46 1510 66
rect 1474 38 1510 46
rect 1616 -28 1631 -19
rect 1002 -43 1631 -28
<< polycont >>
rect 324 153 344 173
rect -104 46 -84 66
rect 541 46 561 66
rect 769 54 789 74
rect 1278 138 1296 156
rect 1482 46 1502 66
<< locali >>
rect -510 231 -504 252
rect -363 236 173 252
rect -486 231 -467 232
rect -363 231 -268 236
rect -249 231 -230 232
rect -127 231 173 236
rect 192 231 211 232
rect 314 231 359 252
rect 377 231 396 232
rect 500 231 1130 252
rect 1136 231 1209 252
rect 1270 231 1316 252
rect 1457 232 1793 252
rect 1334 231 1353 232
rect 1457 231 1811 232
rect 316 173 352 181
rect -109 164 -48 167
rect -109 147 -106 164
rect -89 147 -48 164
rect -109 145 -48 147
rect 316 153 324 173
rect 344 153 352 173
rect 780 154 828 172
rect 1270 156 1304 164
rect 316 145 352 153
rect 127 100 161 104
rect 325 100 342 145
rect 1270 138 1278 156
rect 1296 138 1304 156
rect 1270 133 1304 138
rect 499 110 593 131
rect -561 70 -550 100
rect 293 80 314 87
rect -363 63 -346 78
rect -127 74 -112 80
rect -314 66 -280 70
rect -127 66 -76 74
rect -127 51 -104 66
rect -112 46 -104 51
rect -84 46 -76 66
rect 28 51 145 70
rect 499 68 516 110
rect 761 74 797 82
rect 1066 75 1083 87
rect 1249 79 1270 87
rect 1278 75 1296 133
rect 1436 120 1578 137
rect 1755 93 1773 98
rect 500 63 516 68
rect 533 66 569 74
rect -112 38 -76 46
rect 533 46 541 66
rect 561 46 569 66
rect 761 54 769 74
rect 789 54 797 74
rect 901 58 1083 75
rect 1474 66 1510 74
rect 761 46 797 54
rect 1474 46 1482 66
rect 1502 46 1510 66
rect 1916 63 1931 80
rect 533 38 569 46
rect 1474 38 1510 46
rect -381 -40 -261 -20
rect -145 -40 180 -20
rect 296 -40 366 -20
rect 482 -40 1216 -20
rect 1252 -40 1323 -20
rect 1439 -40 1800 -20
<< viali >>
rect -106 147 -89 164
rect 324 153 344 173
rect 762 154 780 172
rect 1278 138 1296 156
rect -363 78 -346 95
rect -104 46 -84 66
rect 1755 75 1773 93
rect 541 46 561 66
rect 769 54 789 74
rect 1482 46 1502 66
rect 7 2 24 19
rect 656 4 673 21
rect 891 4 908 21
rect 1644 4 1661 21
<< metal1 >>
rect -510 229 -504 252
rect -363 236 173 252
rect -486 231 -467 232
rect -363 229 -268 236
rect -249 231 -230 232
rect -127 229 173 236
rect 192 231 211 232
rect 314 229 359 252
rect 377 231 396 232
rect 500 229 1130 252
rect 1136 229 1209 252
rect 1270 229 1316 252
rect 1457 232 1795 252
rect 1334 231 1353 232
rect 1457 231 1811 232
rect 1457 229 1795 231
rect 316 173 783 181
rect -112 164 -83 171
rect -112 147 -106 164
rect -89 147 -83 164
rect -112 143 -83 147
rect 316 153 324 173
rect 344 172 783 173
rect 344 154 762 172
rect 780 154 783 172
rect 344 153 783 154
rect 316 145 783 153
rect 1267 156 1781 165
rect -112 102 -93 143
rect 1267 138 1278 156
rect 1296 138 1781 156
rect 1267 133 1781 138
rect -369 95 -342 102
rect -140 95 -93 102
rect -369 78 -363 95
rect -346 88 -93 95
rect 1747 93 1781 133
rect -346 78 -126 88
rect -369 77 -126 78
rect -369 72 -342 77
rect 761 74 797 82
rect 1747 75 1755 93
rect 1773 75 1781 93
rect 884 74 924 75
rect -112 66 769 74
rect -112 46 -104 66
rect -84 46 541 66
rect 561 54 769 66
rect 789 66 1510 74
rect 1747 70 1781 75
rect 789 54 1482 66
rect 561 46 1482 54
rect 1502 46 1510 66
rect -112 38 1510 46
rect 1 21 679 24
rect 1 19 656 21
rect 1 2 7 19
rect 24 4 656 19
rect 673 4 679 21
rect 24 2 679 4
rect 1 0 679 2
rect 883 21 1667 24
rect 883 4 891 21
rect 908 4 1644 21
rect 1661 4 1667 21
rect 1 -1 676 0
rect 883 -1 1667 4
rect -381 -45 -261 -15
rect -145 -45 180 -15
rect 296 -45 366 -15
rect 482 -45 1216 -15
rect 1252 -45 1323 -15
rect 1439 -45 1801 -15
use inv1newcell  inv1newcell_0
timestamp 1725972273
transform 1 0 -429 0 1 -28
box -121 -17 66 280
use inv1newcell  inv1newcell_1
timestamp 1725972273
transform 1 0 -193 0 1 -28
box -121 -17 66 280
use inv1newcell  inv1newcell_2
timestamp 1725972273
transform 1 0 248 0 1 -28
box -121 -17 66 280
use inv1newcell  inv1newcell_3
timestamp 1725972273
transform 1 0 434 0 1 -28
box -121 -17 66 280
use inv1newcell  inv1newcell_4
timestamp 1725972273
transform 1 0 1204 0 1 -28
box -121 -17 66 280
use inv1newcell  inv1newcell_5
timestamp 1725972273
transform 1 0 1391 0 1 -28
box -121 -17 66 280
use inv1newcell  inv1newcell_6
timestamp 1725972273
transform 1 0 1868 0 1 -28
box -121 -17 66 280
use Transmissiongate  Transmissiongate_0
timestamp 1726065883
transform -1 0 685 0 1 0
box -82 -19 112 236
use Transmissiongate  Transmissiongate_1
timestamp 1726065883
transform -1 0 920 0 1 0
box -82 -19 112 236
use Transmissiongate  Transmissiongate_2
timestamp 1726065883
transform -1 0 1670 0 1 0
box -82 -19 112 236
use Transmissiongate  Transmissiongate_3
timestamp 1726065883
transform -1 0 36 0 1 0
box -82 -19 112 236
<< labels >>
rlabel locali -556 84 -556 84 7 D
port 1 w
rlabel locali -298 68 -298 68 5 clk
port 2 s
rlabel locali 1929 71 1929 71 7 Q
port 4 w
rlabel metal1 -328 -29 -328 -29 1 gnd
port 6 n
rlabel metal1 -326 242 -326 242 1 vdd
port 5 n
rlabel locali -356 69 -356 69 1 Dbar
rlabel locali -121 63 -121 63 1 clk_inv
rlabel locali 510 77 510 77 1 3
rlabel locali 1077 79 1077 79 1 4
rlabel locali 1266 80 1266 80 1 Qin
rlabel locali 1463 127 1463 127 1 5
rlabel locali 310 80 310 80 1 2
rlabel locali 144 102 144 102 1 1
<< end >>
