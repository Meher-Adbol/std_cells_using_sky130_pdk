module inv1newcell (
    input wire A,
	 output wire Y);

assign Y = ~A;      

endmodule 
