VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFF
  CLASS BLOCK ;
  FOREIGN DFF ;
  ORIGIN 5.610 0.450 ;
  SIZE 24.950 BY 2.970 ;
  PIN D
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT -5.610 0.700 -5.160 1.000 ;
    END
  END D
  PIN clk
    ANTENNAGATEAREA 0.756000 ;
    PORT
      LAYER li1 ;
        RECT -3.140 0.660 -2.800 1.000 ;
    END
  END clk
  PIN Q
    ANTENNADIFFAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 18.890 0.800 19.130 2.140 ;
        RECT 18.890 0.630 19.340 0.800 ;
        RECT 18.890 0.460 19.130 0.630 ;
        RECT 18.870 0.090 19.150 0.460 ;
    END
  END Q
  PIN vdd
    ANTENNADIFFAREA 8.996400 ;
    PORT
      LAYER nwell ;
        RECT -5.100 2.440 19.160 2.520 ;
        RECT -5.100 0.820 19.340 2.440 ;
        RECT -0.760 0.700 1.670 0.820 ;
        RECT 5.730 0.700 10.090 0.820 ;
        RECT 15.580 0.700 17.810 0.820 ;
      LAYER li1 ;
        RECT -5.100 2.320 19.340 2.520 ;
        RECT -5.100 2.310 18.120 2.320 ;
        RECT 18.290 2.310 19.340 2.320 ;
        RECT -4.500 2.140 -4.330 2.310 ;
        RECT -2.140 2.140 -1.970 2.310 ;
        RECT 2.270 2.140 2.440 2.310 ;
        RECT 4.130 2.140 4.300 2.310 ;
        RECT 11.830 2.140 12.000 2.310 ;
        RECT 13.700 2.140 13.870 2.310 ;
        RECT 18.470 2.140 18.640 2.310 ;
        RECT -4.930 1.080 -4.290 2.140 ;
        RECT -2.570 1.080 -1.930 2.140 ;
        RECT 0.550 0.930 0.960 2.120 ;
        RECT 1.840 1.080 2.480 2.140 ;
        RECT 3.700 1.080 4.340 2.140 ;
        RECT 7.040 0.930 7.450 2.120 ;
        RECT 9.390 0.930 9.800 2.120 ;
        RECT 11.400 1.080 12.040 2.140 ;
        RECT 13.270 1.080 13.910 2.140 ;
        RECT 16.890 0.930 17.300 2.120 ;
        RECT 18.040 1.080 18.680 2.140 ;
      LAYER met1 ;
        RECT -5.100 2.290 19.340 2.520 ;
    END
  END vdd
  PIN gnd
    ANTENNADIFFAREA 2.087400 ;
    PORT
      LAYER li1 ;
        RECT -4.940 0.090 -4.270 0.460 ;
        RECT -2.580 0.090 -1.910 0.460 ;
        RECT 1.830 0.090 2.500 0.460 ;
        RECT 3.690 0.090 4.360 0.460 ;
        RECT 11.390 0.090 12.060 0.460 ;
        RECT 13.260 0.090 13.930 0.460 ;
        RECT 18.030 0.090 18.700 0.460 ;
        RECT -4.490 -0.200 -4.320 0.090 ;
        RECT -2.130 -0.200 -1.960 0.090 ;
        RECT 2.280 -0.200 2.450 0.090 ;
        RECT 4.140 -0.200 4.310 0.090 ;
        RECT 11.840 -0.200 12.010 0.090 ;
        RECT 13.710 -0.200 13.880 0.090 ;
        RECT 18.480 -0.200 18.650 0.090 ;
        RECT -4.970 -0.400 19.160 -0.200 ;
      LAYER met1 ;
        RECT -4.970 -0.450 19.160 -0.150 ;
    END
  END gnd
  OBS
      LAYER li1 ;
        RECT -4.080 0.800 -3.840 2.140 ;
        RECT -3.630 0.800 -3.460 0.950 ;
        RECT -4.080 0.630 -3.460 0.800 ;
        RECT -1.720 0.800 -1.480 2.140 ;
        RECT -0.560 1.670 -0.200 2.040 ;
        RECT -1.090 1.450 -0.200 1.670 ;
        RECT -0.560 0.930 -0.200 1.450 ;
        RECT -0.010 0.930 0.370 2.040 ;
        RECT -1.720 0.740 -1.120 0.800 ;
        RECT -1.720 0.630 -0.760 0.740 ;
        RECT -4.080 0.460 -3.840 0.630 ;
        RECT -1.720 0.460 -1.480 0.630 ;
        RECT -1.270 0.510 -0.760 0.630 ;
        RECT -4.100 0.090 -3.820 0.460 ;
        RECT -1.740 0.090 -1.460 0.460 ;
        RECT -1.120 0.380 -0.760 0.510 ;
        RECT -0.490 0.340 -0.270 0.930 ;
        RECT 0.060 0.700 0.280 0.930 ;
        RECT 1.270 0.700 1.610 1.040 ;
        RECT 2.690 0.870 2.930 2.140 ;
        RECT 3.160 1.450 3.520 1.810 ;
        RECT 3.250 1.000 3.420 1.450 ;
        RECT 3.130 0.870 3.470 1.000 ;
        RECT 2.690 0.700 3.470 0.870 ;
        RECT 4.550 0.800 4.790 2.140 ;
        RECT 5.930 1.310 6.290 2.040 ;
        RECT 4.990 1.100 6.290 1.310 ;
        RECT 4.990 0.800 5.160 1.100 ;
        RECT 5.930 0.930 6.290 1.100 ;
        RECT 6.480 0.930 6.860 2.040 ;
        RECT 8.280 1.720 8.640 2.040 ;
        RECT 7.620 1.540 8.640 1.720 ;
        RECT 8.280 0.930 8.640 1.540 ;
        RECT 8.830 0.930 9.210 2.040 ;
        RECT 0.060 0.510 1.450 0.700 ;
        RECT 2.690 0.630 3.140 0.700 ;
        RECT 4.550 0.630 5.160 0.800 ;
        RECT 0.060 0.340 0.280 0.510 ;
        RECT 2.690 0.460 2.930 0.630 ;
        RECT 4.550 0.460 4.790 0.630 ;
        RECT -0.560 0.000 -0.200 0.340 ;
        RECT -0.010 0.000 0.350 0.340 ;
        RECT 0.590 0.000 0.960 0.300 ;
        RECT 2.670 0.090 2.950 0.460 ;
        RECT 4.530 0.090 4.810 0.460 ;
        RECT 5.330 0.380 5.690 0.740 ;
        RECT 6.000 0.340 6.220 0.930 ;
        RECT 6.550 0.340 6.770 0.930 ;
        RECT 7.610 0.460 7.970 0.820 ;
        RECT 8.350 0.340 8.570 0.930 ;
        RECT 8.900 0.750 9.120 0.930 ;
        RECT 10.830 0.870 11.170 1.000 ;
        RECT 10.660 0.750 11.170 0.870 ;
        RECT 8.900 0.700 11.170 0.750 ;
        RECT 12.250 0.870 12.490 2.140 ;
        RECT 12.700 1.330 13.040 1.640 ;
        RECT 14.120 1.370 14.360 2.140 ;
        RECT 15.780 1.370 16.140 2.040 ;
        RECT 12.780 1.000 12.960 1.330 ;
        RECT 14.120 1.200 16.140 1.370 ;
        RECT 12.700 0.870 13.040 1.000 ;
        RECT 12.250 0.700 13.040 0.870 ;
        RECT 14.120 0.800 14.360 1.200 ;
        RECT 15.780 0.930 16.140 1.200 ;
        RECT 16.330 0.930 16.710 2.040 ;
        RECT 8.900 0.580 10.830 0.700 ;
        RECT 12.250 0.630 12.700 0.700 ;
        RECT 14.120 0.630 14.570 0.800 ;
        RECT 8.900 0.340 9.120 0.580 ;
        RECT 12.250 0.460 12.490 0.630 ;
        RECT 14.120 0.460 14.360 0.630 ;
        RECT 5.930 0.000 6.290 0.340 ;
        RECT 6.480 0.000 6.840 0.340 ;
        RECT 7.080 0.000 7.450 0.300 ;
        RECT 8.280 0.000 8.640 0.340 ;
        RECT 8.830 0.000 9.190 0.340 ;
        RECT 9.430 0.000 9.800 0.300 ;
        RECT 12.230 0.090 12.510 0.460 ;
        RECT 14.100 0.090 14.380 0.460 ;
        RECT 14.740 0.380 15.100 0.740 ;
        RECT 15.850 0.340 16.070 0.930 ;
        RECT 16.400 0.340 16.620 0.930 ;
        RECT 17.470 0.700 17.810 1.000 ;
        RECT 15.780 0.000 16.140 0.340 ;
        RECT 16.330 0.000 16.690 0.340 ;
        RECT 16.930 0.000 17.300 0.300 ;
      LAYER met1 ;
        RECT -1.120 1.430 -0.830 1.710 ;
        RECT 3.160 1.450 7.830 1.810 ;
        RECT -1.120 1.020 -0.930 1.430 ;
        RECT 12.670 1.330 17.810 1.650 ;
        RECT -3.690 0.950 -3.420 1.020 ;
        RECT -1.400 0.950 -0.930 1.020 ;
        RECT -3.690 0.880 -0.930 0.950 ;
        RECT -3.690 0.770 -1.260 0.880 ;
        RECT -3.690 0.720 -3.420 0.770 ;
        RECT 7.610 0.740 7.970 0.820 ;
        RECT 8.840 0.740 9.240 0.750 ;
        RECT -1.120 0.380 15.100 0.740 ;
        RECT 17.470 0.700 17.810 1.330 ;
        RECT 0.010 0.000 6.790 0.240 ;
        RECT 0.010 -0.010 6.760 0.000 ;
        RECT 8.830 -0.010 16.670 0.240 ;
  END
END DFF
END LIBRARY

