* Name: Aditya Tare (24M1169), Gautam Govindaraju (24M1166), Ritoo Verma (24M1185), Sachin Soneria (24M1178)
* EE671 - Course Project 01 Group 12
* 3 Input NAND Gate (first input inverted)

*Including sky130 device model
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* Define power supply
Vdd Vdd gnd DC 1.8

* Define input signals
* Vin1 a gnd pulse(0 1.8 42.5ns 20ps 20ps 40ns 80ns)
* Vin2 b gnd pulse(0 1.8 24.5ns 20ps 20ps 20ns 40ns)
* Vin3 c gnd pulse(0 1.8 12.5ns 20ps 20ps 10ns 20ns)
Vin1 a gnd DC 0
Vin2 b gnd DC 1.8
Vin3 c gnd PULSE(0 1.8 0 10ps 10ps 1ns 3ns)

.subckt not1 Vdd vss a z
XM01 z a Vdd Vdd skY130_fd_pr__pfet_01v8 l=0.15 w=1.26 as=0.378 ad=0.378 ps=3.12 pd=3.12
XM02 z a gnd gnd skY130_fd_pr__nfet_01v8 l=0.15 w=0.42 as=0.12 ad=0.12 ps=1.4 pd=1.4
.ends

.subckt nand3 Ain Bin Cin Y Vdd gnd


X0 Abar Ain Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.378 pd=3.12 as=0.3045 ps=2.83 w=1.26 l=0.15
X1 Abar Ain gnd gnd sky130_fd_pr__nfet_01v8 ad=0.126 pd=1.44 as=0.1155 ps=1.18 w=0.42 l=0.15
X2 Y Abar Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.093333 pd=0.911111 as=0.1015 ps=0.943333 w=0.42 l=0.15
X3 2 Cin gnd gnd sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.1155 ps=1.18 w=0.42 l=0.15
X4 4 Bin 3 gnd sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.084 ps=0.82 w=0.42 l=0.15
X5 Y Abar Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.093333 pd=0.911111 as=0.1015 ps=0.943333 w=0.42 l=0.15
X6 Vdd Cin Y Vdd sky130_fd_pr__pfet_01v8 ad=0.1015 pd=0.943333 as=0.093333 ps=0.911111 w=0.42 l=0.15
X7 Y Abar 5 gnd sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.093333 as=0.084 ps=0.82 w=0.42 l=0.15
X8 Vdd Bin Y Vdd sky130_fd_pr__pfet_01v8 ad=0.1015 pd=0.943333 as=0.093333 ps=0.911111 w=0.42 l=0.15
X9 Y Abar 6 gnd sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.093333 as=0.084 ps=0.82 w=0.42 l=0.15
X10 Vdd Bin Y Vdd sky130_fd_pr__pfet_01v8 ad=0.1015 pd=0.943333 as=0.093333 ps=0.911111 w=0.42 l=0.15
X11 gnd Cin 1 gnd sky130_fd_pr__nfet_01v8 ad=0.1155 pd=1.18 as=0.084 ps=0.82 w=0.42 l=0.15
X12 Vdd Abar Y Vdd sky130_fd_pr__pfet_01v8 ad=0.1015 pd=0.943333 as=0.093333 ps=0.911111 w=0.42 l=0.15
X13 3 Bin 2 gnd sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.084 ps=0.82 w=0.42 l=0.15
X14 Y Cin Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.093333 pd=0.911111 as=0.1015 ps=0.943333 w=0.42 l=0.15
X15 5 Bin 4 gnd sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.084 ps=0.82 w=0.42 l=0.15
X16 Y Cin Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.093333 pd=0.911111 as=0.1015 ps=0.943333 w=0.42 l=0.15
X17 6 Abar Y gnd sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.112 ps=1.093333 w=0.42 l=0.15
X18 Y Bin Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.093333 pd=0.911111 as=0.1015 ps=0.943333 w=0.42 l=0.15
X19 1 Cin gnd gnd sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.1155 ps=1.18 w=0.42 l=0.15
C0 gnd 6 0.008175f
C1 Cin Y 0.112245f
C2 Cin 3 5.99e-20
C3 3 Y 0.013389f
C4 gnd 5 0.008119f
C5 Ain Y 6.47e-19
C6 Ain 3 1.37e-20
C7 Cin 4 4.45e-20
C8 gnd Abar 0.028534f
C9 Cin Vdd 0.224506f
C10 Cin Bin 0.151326f
C11 Cin 2 0.00278f
C12 4 Y 0.013535f
C13 Vdd Y 0.714268f
C14 Bin Y 0.10443f
C15 3 4 0.022948f
C16 2 Y 0.013316f
C17 3 Vdd 0.001508f
C18 Ain 4 1.81e-20
C19 Ain Vdd 0.120775f
C20 3 Bin 0.00917f
C21 2 3 0.023542f
C22 Ain Bin 1.09e-19
C23 Ain 2 1.07e-20
C24 Cin 6 2.05e-21
C25 4 Vdd 7.46e-19
C26 gnd 1 0.008067f
C27 4 Bin 0.009169f
C28 Bin Vdd 0.475151f
C29 6 Y 0.061468f
C30 2 Vdd 7.46e-19
C31 2 Bin 0.002909f
C32 6 Ain 5.76e-20
C33 Cin 5 3.44e-20
C34 6 Vdd 0.001508f
C35 Y 5 0.037969f
C36 Cin Abar 5.77e-20
C37 Ain 5 2.5e-20
C38 Y Abar 0.171193f
C39 Ain Abar 0.046385f
C40 4 5 0.023542f
C41 Vdd 5 0.001508f
C42 Bin 5 0.002677f
C43 Vdd Abar 0.396396f
C44 Cin 1 0.009377f
C45 gnd Cin 0.026634f
C46 Bin Abar 0.052035f
C47 1 Y 0.013255f
C48 gnd Y 0.043914f
C49 gnd 3 0.008097f
C50 1 Ain 7.1e-21
C51 gnd Ain 9.68e-21
C52 6 Abar 0.00917f
C53 gnd 4 0.008106f
C54 1 Vdd 7.46e-19
C55 gnd Vdd 0.15604f
C56 gnd Bin 0.020086f
C57 gnd 2 0.008091f
C58 5 Abar 0.002712f
C59 gnd 0 0.560006f
C60 Y 0 0.35291f
C61 Cin 0 0.666468f
C62 Bin 0 0.790311f
C63 6 0 0.034171f
C64 5 0 0.034681f
C65 4 0 0.034306f
C66 3 0 0.034452f
C67 2 0 0.058699f
C68 1 0 0.082385f
C69 Abar 0 0.716198f
C70 Ain 0 0.318198f
C71 Vdd 0 2.065253f

.ends

Xnand1 a b c out Vdd gnd nand3
*Xnot1 Vdd gnd out InvertedOut not1
Cload out gnd 0.5f

* Define simulation Control
.tran 0.1ps 20ns 0 1p

.control

* run
* plot V(out) V(a)+2
* let StaticPower = I(Vdd) * Vdd
* print StaticPower



******************** DYNAMIC POWER CHARACTERISTICS ********************

foreach val 0.5e-15 10e-15 100e-15
	foreach varx 10e-12 100e-12 1000e-12
		let a1=0
		let a2=$varx
		let b1=(3000e-12 - $varx)
		let b2=(3000e-12)
		let hold=(3000e-12 - 2 * $varx)
        alter @Cload $val
		alter @Vin3[PULSE] [ 0 1.8 0 $varx $varx $&hold 6n ]
		echo CLoad is $val InputSlew is $varx
		echo rise from 0 to $&a2
		echo fall from $&b1 to $&b2
		run	
		meas tran Ipeak_rise MAX I(Vdd) from=0 to=$&a2
		meas tran Ipeak_fall MIN I(Vdd) from=$&b1 to=$&b2
		let RISE_POWER= (0.5* $varx * Ipeak_rise *1.8)/$&b2
		let FALL_POWER= (0.5 *$varx * Ipeak_fall * 1.8)/$&b2
		print RISE_POWER
		print FALL_POWER
		reset
	end	
end



******************** TIMING CHARACTERISTICS ********************

* foreach val 0.5e-15 10e-15 100e-15
	* foreach varx 10e-12 100e-12 1000e-12
        * alter @Cload $val
		* alter @Vin3[PULSE] [ 0 1.8 0 $varx $varx 4n 10n ]
		* echo CLoad is $val InputSlew is $varx
		* run
		* meas tran T_RISE TRIG v(out) VAL = 0.36 RISE = 1 TARG v(out) VAL = 1.44 RISE = 1
		* meas tran T_FALL TRIG v(out) VAL = 1.44 FALL = 1 TARG v(out) VAL = 0.36 FALL = 1
		* meas tran CELL_RISE_DELAY TRIG v(c)  VAL = 0.9 FALL = 1 TARG v(out) VAL = 0.9 RISE = 1
		* meas tran CELL_FALL_DELAY TRIG v(c)  VAL = 0.9 RISE = 1 TARG v(out) VAL = 0.9 FALL = 1	
		* plot V(out) V(c)+2
		* reset
	* end	
* end

******************** INPUT CAPACITANCE ********************
* In this part we first inject a known voltage source and we integrate the current during falling and rising edges of the voltage source , these values
* of current are used to calculate input capacitance.
* meas tran AI_integ_rise INTEG I(Vin1) from=0p to =500p
* meas tran AI_integ_fall INTEG I(Vin1) from=1500p to =2000p
* let AInputCapRise=AI_integ_rise/1.8
* let AInputCapFall=AI_integ_fall/1.8
* let AAvg_Cap=(AInputCapRise+AInputCapFall)/2
* print AInputCapRise AInputCapFall AAvg_Cap

* meas tran BI_integ_rise INTEG I(Vin2) from=0p to =500p
* meas tran BI_integ_fall INTEG I(Vin2) from=1500p to =2000p
* let BInputCapRise=BI_integ_rise/1.8
* let BInputCapFall=BI_integ_fall/1.8
* let BAvg_Cap=(BInputCapRise+BInputCapFall)/2
* print BInputCapRise BInputCapFall BAvg_Cap

* meas tran CI_integ_rise INTEG I(Vin3) from=0p to =500p
* meas tran CI_integ_fall INTEG I(Vin3) from=1500p to =2000p
* let CInputCapRise=CI_integ_rise/1.8
* let CInputCapFall=CI_integ_fall/1.8
* let CAvg_Cap=(CInputCapRise+CInputCapFall)/2
* print CInputCapRise CInputCapFall CAvg_Cap

set color0=white
set color1=black
set color2=blue
set color3=green
set color4=red
set color5=purple
set xbrushwidth=4

.endc
