module buff(input a,
	    output y);
	    
assign y=a;
endmodule
