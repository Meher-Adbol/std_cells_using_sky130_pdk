magic
tech sky130A
timestamp 1726413032
<< nwell >>
rect -55 1356 213 1519
rect 344 1357 603 1583
<< nmos >>
rect 105 1254 120 1296
rect 540 1186 555 1246
<< pmos >>
rect 105 1374 120 1501
rect 540 1375 555 1565
<< ndiff >>
rect 75 1284 105 1296
rect 75 1264 81 1284
rect 98 1264 105 1284
rect 75 1254 105 1264
rect 120 1284 150 1296
rect 120 1264 128 1284
rect 145 1264 150 1284
rect 120 1254 150 1264
rect 510 1235 540 1246
rect 510 1194 517 1235
rect 534 1194 540 1235
rect 510 1186 540 1194
rect 555 1235 585 1246
rect 555 1194 562 1235
rect 579 1194 585 1235
rect 555 1186 585 1194
<< pdiff >>
rect 75 1486 105 1501
rect 75 1386 81 1486
rect 99 1386 105 1486
rect 75 1374 105 1386
rect 120 1486 150 1501
rect 120 1386 126 1486
rect 144 1386 150 1486
rect 120 1374 150 1386
rect 510 1552 540 1565
rect 510 1390 516 1552
rect 533 1390 540 1552
rect 510 1375 540 1390
rect 555 1552 585 1565
rect 555 1390 562 1552
rect 579 1390 585 1552
rect 555 1375 585 1390
<< ndiffc >>
rect 81 1264 98 1284
rect 128 1264 145 1284
rect 517 1194 534 1235
rect 562 1194 579 1235
<< pdiffc >>
rect 81 1386 99 1486
rect 126 1386 144 1486
rect 516 1390 533 1552
rect 562 1390 579 1552
<< psubdiff >>
rect 32 1285 75 1296
rect 32 1265 44 1285
rect 61 1265 75 1285
rect 32 1254 75 1265
rect 460 1234 510 1246
rect 460 1193 477 1234
rect 494 1193 510 1234
rect 460 1186 510 1193
<< nsubdiff >>
rect 365 1549 440 1565
rect -30 1484 45 1501
rect -30 1391 -14 1484
rect 25 1391 45 1484
rect -30 1374 45 1391
rect 365 1385 384 1549
rect 420 1385 440 1549
rect 365 1375 440 1385
<< psubdiffcont >>
rect 44 1265 61 1285
rect 477 1193 494 1234
<< nsubdiffcont >>
rect -14 1391 25 1484
rect 384 1385 420 1549
<< poly >>
rect 540 1565 555 1583
rect 105 1501 120 1514
rect -100 1345 -60 1355
rect 105 1345 120 1374
rect -100 1325 -90 1345
rect -70 1328 120 1345
rect -70 1325 -60 1328
rect -100 1315 -60 1325
rect 105 1296 120 1328
rect 290 1334 333 1337
rect 540 1334 555 1375
rect 290 1327 555 1334
rect 290 1307 301 1327
rect 321 1307 555 1327
rect 290 1304 555 1307
rect 290 1297 333 1304
rect 105 1230 120 1254
rect 540 1246 555 1304
rect 540 1172 555 1186
<< polycont >>
rect -90 1325 -70 1345
rect 301 1307 321 1327
<< locali >>
rect -15 1685 27 1690
rect -15 1665 -5 1685
rect 15 1665 27 1685
rect -15 1501 27 1665
rect 384 1684 418 1689
rect 384 1664 391 1684
rect 411 1664 418 1684
rect 384 1565 418 1664
rect 365 1552 538 1565
rect 365 1549 516 1552
rect -30 1486 105 1501
rect -30 1484 81 1486
rect -30 1391 -14 1484
rect 25 1391 81 1484
rect -30 1386 81 1391
rect 99 1386 105 1486
rect -30 1374 105 1386
rect 122 1486 149 1500
rect 122 1386 126 1486
rect 144 1386 149 1486
rect 122 1376 149 1386
rect -100 1345 -60 1355
rect -100 1325 -90 1345
rect -70 1325 -60 1345
rect -100 1315 -60 1325
rect 131 1331 149 1376
rect 365 1385 384 1549
rect 420 1390 516 1549
rect 533 1390 538 1552
rect 420 1385 538 1390
rect 365 1375 538 1385
rect 555 1552 585 1565
rect 555 1390 562 1552
rect 579 1390 585 1552
rect 555 1375 585 1390
rect 562 1346 585 1375
rect 290 1331 333 1337
rect 131 1327 333 1331
rect 131 1307 301 1327
rect 321 1307 333 1327
rect 131 1306 333 1307
rect 131 1296 149 1306
rect 290 1297 333 1306
rect 562 1321 725 1346
rect 32 1285 105 1296
rect 32 1265 44 1285
rect 61 1284 105 1285
rect 61 1265 81 1284
rect 32 1264 81 1265
rect 98 1264 105 1284
rect 32 1254 105 1264
rect 122 1284 149 1296
rect 122 1264 128 1284
rect 145 1264 149 1284
rect 122 1254 149 1264
rect 34 1140 68 1254
rect 562 1246 585 1321
rect 460 1235 537 1246
rect 460 1234 517 1235
rect 460 1193 477 1234
rect 494 1194 517 1234
rect 534 1194 537 1235
rect 494 1193 537 1194
rect 460 1186 537 1193
rect 555 1235 585 1246
rect 555 1194 562 1235
rect 579 1194 585 1235
rect 555 1186 585 1194
rect 34 1120 40 1140
rect 60 1120 68 1140
rect 34 1115 68 1120
rect 466 1140 501 1186
rect 466 1120 473 1140
rect 493 1120 501 1140
rect 466 1115 501 1120
<< viali >>
rect -5 1665 15 1685
rect 391 1664 411 1684
rect 40 1120 60 1140
rect 473 1120 493 1140
<< metal1 >>
rect -105 1685 734 1690
rect -105 1665 -5 1685
rect 15 1684 734 1685
rect 15 1665 391 1684
rect -105 1664 391 1665
rect 411 1664 734 1684
rect -105 1659 734 1664
rect -85 1140 705 1145
rect -85 1120 40 1140
rect 60 1120 473 1140
rect 493 1120 705 1140
rect -85 1115 705 1120
<< labels >>
rlabel metal1 -85 1130 -85 1130 7 Vss
port 3 w
rlabel metal1 -105 1674 -105 1674 7 Vdd
port 2 w
rlabel locali 725 1335 725 1335 3 out2
port 4 e
rlabel locali -100 1335 -100 1335 7 in
port 1 w
<< end >>
