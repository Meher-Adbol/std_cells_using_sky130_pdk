magic
tech sky130A
timestamp 1726067859
<< nwell >>
rect -551 182 191 266
<< nmos >>
rect -445 64 -430 106
rect -390 64 -375 106
rect -335 64 -320 106
rect -280 64 -265 106
rect -225 64 -210 106
rect -170 64 -155 106
rect -115 64 -100 106
rect -60 64 -45 106
rect -5 64 10 106
<< pmos >>
rect -445 200 -430 242
rect -390 200 -375 242
rect -335 200 -320 242
rect -280 200 -265 242
rect -225 200 -210 242
rect -170 200 -155 242
rect -115 200 -100 242
rect -60 200 -45 242
rect -5 200 10 242
<< ndiff >>
rect -485 100 -445 106
rect -485 70 -475 100
rect -455 70 -445 100
rect -485 64 -445 70
rect -430 100 -390 106
rect -430 70 -420 100
rect -400 70 -390 100
rect -430 64 -390 70
rect -375 100 -335 106
rect -375 70 -365 100
rect -345 70 -335 100
rect -375 64 -335 70
rect -320 100 -280 106
rect -320 70 -310 100
rect -290 70 -280 100
rect -320 64 -280 70
rect -265 100 -225 106
rect -265 70 -255 100
rect -235 70 -225 100
rect -265 64 -225 70
rect -210 100 -170 106
rect -210 70 -199 100
rect -179 70 -170 100
rect -210 64 -170 70
rect -155 100 -115 106
rect -155 70 -144 100
rect -124 70 -115 100
rect -155 64 -115 70
rect -100 100 -60 106
rect -100 70 -89 100
rect -69 70 -60 100
rect -100 64 -60 70
rect -45 100 -5 106
rect -45 70 -35 100
rect -15 70 -5 100
rect -45 64 -5 70
rect 10 100 50 106
rect 10 70 20 100
rect 40 70 50 100
rect 10 64 50 70
<< pdiff >>
rect -485 236 -445 242
rect -485 206 -475 236
rect -455 206 -445 236
rect -485 200 -445 206
rect -430 236 -390 242
rect -430 206 -420 236
rect -400 206 -390 236
rect -430 200 -390 206
rect -375 236 -335 242
rect -375 206 -365 236
rect -345 206 -335 236
rect -375 200 -335 206
rect -320 236 -280 242
rect -320 206 -310 236
rect -290 206 -280 236
rect -320 200 -280 206
rect -265 236 -225 242
rect -265 206 -255 236
rect -235 206 -225 236
rect -265 200 -225 206
rect -210 236 -170 242
rect -210 206 -200 236
rect -180 206 -170 236
rect -210 200 -170 206
rect -155 236 -115 242
rect -155 206 -145 236
rect -125 206 -115 236
rect -155 200 -115 206
rect -100 236 -60 242
rect -100 206 -90 236
rect -70 206 -60 236
rect -100 200 -60 206
rect -45 236 -5 242
rect -45 206 -35 236
rect -15 206 -5 236
rect -45 200 -5 206
rect 10 236 50 242
rect 10 206 20 236
rect 40 206 50 236
rect 10 200 50 206
<< ndiffc >>
rect -475 70 -455 100
rect -420 70 -400 100
rect -365 70 -345 100
rect -310 70 -290 100
rect -255 70 -235 100
rect -199 70 -179 100
rect -144 70 -124 100
rect -89 70 -69 100
rect -35 70 -15 100
rect 20 70 40 100
<< pdiffc >>
rect -475 206 -455 236
rect -420 206 -400 236
rect -365 206 -345 236
rect -310 206 -290 236
rect -255 206 -235 236
rect -200 206 -180 236
rect -145 206 -125 236
rect -90 206 -70 236
rect -35 206 -15 236
rect 20 206 40 236
<< psubdiff >>
rect 50 100 93 106
rect 50 70 60 100
rect 81 70 93 100
rect 50 64 93 70
<< nsubdiff >>
rect 50 236 93 242
rect 50 206 60 236
rect 81 206 93 236
rect 50 200 93 206
<< psubdiffcont >>
rect 60 70 81 100
<< nsubdiffcont >>
rect 60 206 81 236
<< poly >>
rect -541 286 -265 301
rect -541 250 -526 286
rect -552 242 -516 250
rect -445 242 -430 257
rect -390 250 -320 265
rect -390 242 -375 250
rect -335 242 -320 250
rect -280 242 -265 286
rect -225 250 -155 265
rect -225 242 -210 250
rect -170 242 -155 250
rect -115 250 -45 265
rect -115 242 -100 250
rect -60 242 -45 250
rect -5 242 10 255
rect -552 222 -544 242
rect -524 222 -516 242
rect -552 214 -516 222
rect -445 192 -430 200
rect -390 192 -375 200
rect -445 177 -375 192
rect -536 129 -500 134
rect -536 126 -375 129
rect -536 106 -528 126
rect -508 114 -375 126
rect -508 106 -500 114
rect -445 106 -430 114
rect -390 106 -375 114
rect -335 106 -320 200
rect -280 192 -265 200
rect -225 192 -210 200
rect -280 177 -210 192
rect -280 114 -210 129
rect -280 106 -265 114
rect -225 106 -210 114
rect -170 106 -155 200
rect -115 106 -100 200
rect -60 192 -45 200
rect -5 192 10 200
rect -60 177 10 192
rect 93 151 129 159
rect 93 138 101 151
rect 63 131 101 138
rect 121 131 129 151
rect 63 129 129 131
rect -60 123 129 129
rect -60 114 78 123
rect -60 106 -45 114
rect -5 106 10 114
rect -536 98 -500 106
rect -445 51 -430 64
rect -390 56 -375 64
rect -335 56 -320 64
rect -390 41 -320 56
rect -280 51 -265 64
rect -225 56 -210 64
rect -170 56 -155 64
rect -225 41 -155 56
rect -115 56 -100 64
rect -60 56 -45 64
rect -115 41 -45 56
rect -5 51 10 64
<< polycont >>
rect -544 222 -524 242
rect -528 106 -508 126
rect 101 131 121 151
<< locali >>
rect -695 303 -691 323
rect -630 321 319 324
rect -630 304 -419 321
rect -401 304 22 321
rect 39 304 319 321
rect -630 303 319 304
rect -552 242 -516 250
rect -419 242 -401 303
rect -309 244 -291 303
rect -253 266 -16 283
rect -552 222 -544 242
rect -524 222 -516 242
rect -552 214 -516 222
rect -483 236 -446 242
rect -483 206 -475 236
rect -455 206 -446 236
rect -483 203 -446 206
rect -428 236 -392 242
rect -428 206 -420 236
rect -400 206 -392 236
rect -428 203 -392 206
rect -373 236 -337 242
rect -373 206 -365 236
rect -345 206 -337 236
rect -373 203 -337 206
rect -318 236 -282 244
rect -253 242 -236 266
rect -144 242 -126 266
rect -34 242 -16 266
rect 21 242 39 303
rect -318 206 -310 236
rect -290 206 -282 236
rect -318 203 -282 206
rect -263 236 -227 242
rect -263 206 -255 236
rect -235 206 -227 236
rect -263 203 -227 206
rect -208 236 -172 242
rect -208 206 -200 236
rect -180 206 -172 236
rect -208 203 -172 206
rect -153 236 -117 242
rect -153 206 -145 236
rect -125 206 -117 236
rect -153 203 -117 206
rect -98 236 -62 242
rect -98 206 -90 236
rect -70 206 -62 236
rect -98 203 -62 206
rect -43 236 -7 242
rect -43 206 -35 236
rect -15 206 -7 236
rect -43 203 -7 206
rect 12 236 90 242
rect 12 206 20 236
rect 40 206 60 236
rect 81 206 90 236
rect 12 203 90 206
rect -748 142 -737 172
rect -551 135 -519 152
rect -536 134 -519 135
rect -474 141 -456 203
rect -364 141 -346 203
rect -309 176 -291 203
rect -199 176 -181 203
rect -309 158 -199 176
rect -144 141 -126 203
rect -89 176 -71 203
rect 20 176 40 203
rect -71 158 40 176
rect -474 137 -126 141
rect -536 126 -500 134
rect -536 106 -528 126
rect -508 106 -500 126
rect -536 98 -500 106
rect -474 124 -144 137
rect -474 100 -456 124
rect -364 100 -346 124
rect -146 120 -144 124
rect -127 120 -126 137
rect 93 151 129 159
rect 93 131 101 151
rect 121 131 129 151
rect 337 135 362 152
rect 93 123 129 131
rect -146 118 -126 120
rect -483 70 -475 100
rect -455 70 -447 100
rect -428 70 -420 100
rect -400 70 -392 100
rect -373 70 -365 100
rect -345 70 -337 100
rect -318 70 -310 100
rect -290 70 -282 100
rect -263 70 -255 100
rect -235 70 -227 100
rect -207 70 -199 100
rect -179 70 -171 100
rect -152 70 -144 100
rect -124 70 -116 100
rect -97 70 -89 100
rect -69 70 -61 100
rect -43 70 -35 100
rect -15 70 -7 100
rect 12 70 20 100
rect 40 70 60 100
rect 81 70 89 100
rect -88 52 -70 70
rect 21 69 89 70
rect 21 52 39 69
rect -694 32 -683 52
rect -568 35 22 52
rect 39 35 203 52
rect -568 32 203 35
rect 319 32 365 52
<< viali >>
rect -419 304 -401 321
rect 22 304 39 321
rect -199 158 -181 176
rect -89 158 -71 176
rect -144 120 -127 137
rect 158 147 176 165
rect 22 35 39 52
<< metal1 >>
rect -695 324 365 330
rect -695 301 -691 324
rect -630 321 365 324
rect -630 304 -419 321
rect -401 304 22 321
rect 39 304 365 321
rect -630 301 365 304
rect -695 298 365 301
rect -311 176 -289 298
rect -204 176 -175 179
rect -311 158 -199 176
rect -181 158 -175 176
rect -204 155 -175 158
rect -95 176 -66 179
rect 18 176 42 298
rect -95 158 -89 176
rect -71 158 42 176
rect 150 165 184 172
rect -95 155 -66 158
rect 150 147 158 165
rect 176 147 184 165
rect 150 140 184 147
rect -150 137 184 140
rect -150 120 -144 137
rect -127 120 184 137
rect -150 116 184 120
rect -695 52 -684 57
rect -568 52 203 57
rect -695 32 -683 52
rect -568 35 22 52
rect 39 35 203 52
rect -695 27 -684 32
rect -568 27 203 35
rect 319 27 365 57
use inv1newcell  inv1newcell_0 /mnt/c/WINDOWS/system32/new_pdk_sky/layout/course_project
timestamp 1725972273
transform 1 0 -616 0 1 44
box -121 -17 66 280
use inv1newcell  inv1newcell_1
timestamp 1725972273
transform 1 0 271 0 1 44
box -121 -17 66 280
<< labels >>
rlabel locali -544 232 -544 232 7 Bin
port 5 w
rlabel locali 101 141 101 141 7 Cin
port 6 w
rlabel metal1 -144 128 -144 128 7 Y
port 7 w
rlabel locali 359 143 359 143 7 Ybar
port 8 w
rlabel space -673 312 -673 312 7 Vdd
port 2 w
rlabel space -672 44 -672 44 7 gnd
port 3 w
rlabel locali -550 143 -550 143 3 Abar
port 4 e
rlabel locali -746 156 -746 156 3 Ain
port 1 e
<< end >>
