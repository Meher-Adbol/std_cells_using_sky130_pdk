magic
tech sky130A
timestamp 1726412341
<< nwell >>
rect -147 72 38 235
rect 167 92 388 255
rect 663 72 848 235
rect -147 71 -25 72
rect 663 71 785 72
<< nmos >>
rect -25 -5 -10 37
rect 280 15 295 57
rect 325 15 340 57
rect 470 15 485 57
rect 515 15 530 57
rect 785 -5 800 37
<< pmos >>
rect -25 90 -10 217
rect 280 110 295 237
rect 325 110 340 237
rect 785 90 800 217
<< ndiff >>
rect -55 26 -25 37
rect -55 5 -48 26
rect -31 5 -25 26
rect -55 -5 -25 5
rect -10 26 20 37
rect -10 5 -4 26
rect 13 5 20 26
rect 250 43 280 57
rect 250 25 255 43
rect 273 25 280 43
rect 250 15 280 25
rect 295 43 325 57
rect 295 25 301 43
rect 319 25 325 43
rect 295 15 325 25
rect 340 43 370 57
rect 340 25 347 43
rect 365 25 370 43
rect 340 15 370 25
rect 440 43 470 57
rect 440 25 445 43
rect 463 25 470 43
rect 440 15 470 25
rect 485 43 515 57
rect 485 25 491 43
rect 509 25 515 43
rect 485 15 515 25
rect 530 43 560 57
rect 530 25 537 43
rect 555 25 560 43
rect 530 15 560 25
rect -10 -5 20 5
rect 755 26 785 37
rect 755 5 762 26
rect 779 5 785 26
rect 755 -5 785 5
rect 800 26 830 37
rect 800 5 806 26
rect 823 5 830 26
rect 800 -5 830 5
<< pdiff >>
rect -55 146 -25 217
rect -55 111 -50 146
rect -33 111 -25 146
rect -55 90 -25 111
rect -10 146 20 217
rect -10 111 -2 146
rect 15 111 20 146
rect -10 90 20 111
rect 250 192 280 237
rect 250 165 255 192
rect 273 165 280 192
rect 250 110 280 165
rect 295 192 325 237
rect 295 165 301 192
rect 319 165 325 192
rect 295 110 325 165
rect 340 192 370 237
rect 340 165 347 192
rect 365 165 370 192
rect 340 110 370 165
rect 755 146 785 217
rect 755 111 760 146
rect 777 111 785 146
rect 755 90 785 111
rect 800 146 830 217
rect 800 111 808 146
rect 825 111 830 146
rect 800 90 830 111
<< ndiffc >>
rect -48 5 -31 26
rect -4 5 13 26
rect 255 25 273 43
rect 301 25 319 43
rect 347 25 365 43
rect 445 25 463 43
rect 491 25 509 43
rect 537 25 555 43
rect 762 5 779 26
rect 806 5 823 26
<< pdiffc >>
rect -50 111 -33 146
rect -2 111 15 146
rect 255 165 273 192
rect 301 165 319 192
rect 347 165 365 192
rect 760 111 777 146
rect 808 111 825 146
<< psubdiff >>
rect 210 44 250 57
rect -95 27 -55 37
rect -95 7 -83 27
rect -66 7 -55 27
rect -95 -5 -55 7
rect 210 27 221 44
rect 238 27 250 44
rect 210 15 250 27
rect 560 44 600 57
rect 560 27 572 44
rect 589 27 600 44
rect 560 15 600 27
rect 715 27 755 37
rect 715 7 727 27
rect 744 7 755 27
rect 715 -5 755 7
<< nsubdiff >>
rect -129 145 -94 217
rect -129 110 -121 145
rect -104 110 -94 145
rect -129 90 -94 110
rect 185 187 215 237
rect 185 160 191 187
rect 209 160 215 187
rect 185 110 215 160
rect 681 145 716 217
rect 681 110 689 145
rect 706 110 716 145
rect 681 90 716 110
<< psubdiffcont >>
rect -83 7 -66 27
rect 221 27 238 44
rect 572 27 589 44
rect 727 7 744 27
<< nsubdiffcont >>
rect -121 110 -104 145
rect 191 160 209 187
rect 689 110 706 145
<< poly >>
rect 280 237 295 250
rect 325 237 340 250
rect -25 217 -10 230
rect 785 217 800 230
rect 445 161 485 170
rect 445 140 453 161
rect 475 160 485 161
rect 475 140 640 160
rect 445 132 485 140
rect 280 92 295 110
rect -25 37 -10 90
rect 65 74 100 82
rect 65 72 73 74
rect 64 55 73 72
rect 65 53 73 55
rect 92 72 100 74
rect 143 75 295 92
rect 143 72 161 75
rect 92 55 161 72
rect 280 57 295 75
rect 325 57 340 110
rect 460 102 494 110
rect 460 83 468 102
rect 486 83 494 102
rect 460 75 494 83
rect 470 57 485 75
rect 515 57 530 80
rect 625 60 640 140
rect 785 60 800 90
rect 92 53 100 55
rect 65 45 100 53
rect 625 45 800 60
rect 785 37 800 45
rect -25 -18 -10 -5
rect 280 -10 295 15
rect 325 -10 340 15
rect 470 -10 485 15
rect 515 -10 530 15
rect 785 -18 800 -5
<< polycont >>
rect 453 140 475 161
rect 73 53 92 74
rect 468 83 486 102
<< locali >>
rect -129 262 -94 267
rect -129 241 -125 262
rect -99 241 -94 262
rect -129 217 -94 241
rect 185 262 215 267
rect 185 242 189 262
rect 210 242 215 262
rect 185 237 215 242
rect 342 263 370 267
rect 342 243 346 263
rect 367 243 370 263
rect -129 146 -27 217
rect -129 145 -50 146
rect -129 110 -121 145
rect -104 111 -50 145
rect -33 111 -27 146
rect -104 110 -27 111
rect -129 90 -27 110
rect -8 146 20 217
rect -8 111 -2 146
rect 15 111 20 146
rect -8 90 20 111
rect 185 192 278 237
rect 185 187 255 192
rect 185 160 191 187
rect 209 165 255 187
rect 273 165 278 192
rect 209 160 278 165
rect 185 110 278 160
rect 297 192 323 237
rect 297 165 301 192
rect 319 165 323 192
rect 297 139 323 165
rect 297 122 302 139
rect 319 122 323 139
rect 297 110 323 122
rect 342 192 370 243
rect 342 165 347 192
rect 365 165 370 192
rect 681 262 716 267
rect 681 242 687 262
rect 708 242 716 262
rect 681 217 716 242
rect 342 110 370 165
rect 395 163 485 170
rect 395 136 401 163
rect 419 161 485 163
rect 419 140 453 161
rect 475 140 485 161
rect 419 136 485 140
rect 395 130 485 136
rect 681 146 783 217
rect 681 145 760 146
rect 681 110 689 145
rect 706 111 760 145
rect 777 111 783 146
rect 706 110 783 111
rect 460 102 494 110
rect 460 92 468 102
rect 0 72 20 90
rect 143 83 468 92
rect 486 83 494 102
rect 681 90 783 110
rect 802 146 830 217
rect 802 111 808 146
rect 825 111 830 146
rect 802 90 830 111
rect 65 74 100 82
rect 65 72 73 74
rect 0 55 73 72
rect 0 37 20 55
rect 65 53 73 55
rect 92 72 100 74
rect 143 75 494 83
rect 143 72 161 75
rect 92 55 161 72
rect 810 72 830 90
rect 92 53 100 55
rect 65 45 100 53
rect -95 27 -27 37
rect -95 7 -83 27
rect -66 26 -27 27
rect -66 7 -48 26
rect -95 5 -48 7
rect -31 5 -27 26
rect -95 -5 -27 5
rect -8 26 20 37
rect -8 5 -4 26
rect 13 5 20 26
rect -8 -5 20 5
rect 210 44 278 57
rect 210 27 221 44
rect 238 43 278 44
rect 238 27 255 43
rect 210 25 255 27
rect 273 25 278 43
rect 210 15 278 25
rect 297 43 323 57
rect 297 25 301 43
rect 319 25 323 43
rect 297 15 323 25
rect 342 51 468 57
rect 342 43 389 51
rect 342 25 347 43
rect 365 25 389 43
rect 415 43 468 51
rect 415 25 445 43
rect 463 25 468 43
rect 342 15 468 25
rect 487 43 513 57
rect 487 25 491 43
rect 509 25 513 43
rect 487 15 513 25
rect 532 44 600 57
rect 532 43 572 44
rect 532 25 537 43
rect 555 27 572 43
rect 589 27 600 44
rect 810 55 848 72
rect 810 37 830 55
rect 555 25 600 27
rect 532 15 600 25
rect -95 -11 -55 -5
rect -95 -28 -88 -11
rect -62 -28 -55 -11
rect -95 -35 -55 -28
rect 210 -11 250 15
rect 210 -28 217 -11
rect 244 -28 250 -11
rect 210 -35 250 -28
rect 300 -15 320 15
rect 490 -15 510 15
rect 300 -35 510 -15
rect 560 -11 600 15
rect 560 -28 567 -11
rect 594 -28 600 -11
rect 560 -35 600 -28
rect 715 27 783 37
rect 715 7 727 27
rect 744 26 783 27
rect 744 7 762 26
rect 715 5 762 7
rect 779 5 783 26
rect 715 -5 783 5
rect 802 26 830 37
rect 802 5 806 26
rect 823 5 830 26
rect 802 -5 830 5
rect 715 -11 755 -5
rect 715 -28 722 -11
rect 748 -28 755 -11
rect 715 -35 755 -28
<< viali >>
rect -125 241 -99 262
rect 189 242 210 262
rect 346 243 367 263
rect 302 122 319 139
rect 687 242 708 262
rect 401 136 419 163
rect 389 25 415 51
rect -88 -28 -62 -11
rect 217 -28 244 -11
rect 567 -28 594 -11
rect 722 -28 748 -11
<< metal1 >>
rect -175 263 848 267
rect -175 262 346 263
rect -175 241 -125 262
rect -99 242 189 262
rect 210 243 346 262
rect 367 262 848 263
rect 367 243 687 262
rect 210 242 687 243
rect 708 242 848 262
rect -99 241 848 242
rect -175 237 848 241
rect 395 163 425 170
rect 395 145 401 163
rect 295 139 401 145
rect 295 122 302 139
rect 319 136 401 139
rect 419 136 425 163
rect 319 130 425 136
rect 319 122 420 130
rect 295 115 420 122
rect 385 51 420 115
rect 385 25 389 51
rect 415 25 420 51
rect 385 15 420 25
rect -175 -11 848 -5
rect -175 -28 -88 -11
rect -62 -28 217 -11
rect 244 -28 567 -11
rect 594 -28 722 -11
rect 748 -28 848 -11
rect -175 -35 848 -28
<< labels >>
rlabel locali 82 82 82 82 7 out
<< end >>
