VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO InverterCell
  CLASS BLOCK ;
  FOREIGN InverterCell ;
  ORIGIN 1.210 0.170 ;
  SIZE 1.870 BY 2.970 ;
  PIN vdd
    ANTENNADIFFAREA 0.831600 ;
    PORT
      LAYER nwell ;
        RECT -0.810 0.980 0.660 2.600 ;
      LAYER li1 ;
        RECT -0.750 2.590 0.660 2.800 ;
        RECT -0.560 2.350 -0.390 2.590 ;
        RECT -0.610 1.240 0.000 2.350 ;
      LAYER met1 ;
        RECT -0.750 2.570 0.660 2.800 ;
    END
  END vdd
  PIN vss
    ANTENNADIFFAREA 0.298200 ;
    PORT
      LAYER li1 ;
        RECT -0.650 0.250 0.020 0.620 ;
        RECT -0.560 0.080 -0.380 0.250 ;
        RECT -0.680 -0.120 0.480 0.080 ;
      LAYER met1 ;
        RECT -0.680 -0.170 0.480 0.130 ;
    END
  END vss
  PIN a
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT -1.210 0.760 -0.870 1.060 ;
    END
  END a
  PIN z
    ANTENNADIFFAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.210 0.960 0.450 2.350 ;
        RECT 0.210 0.790 0.660 0.960 ;
        RECT 0.210 0.620 0.450 0.790 ;
        RECT 0.190 0.250 0.470 0.620 ;
    END
  END z
END InverterCell
END LIBRARY

