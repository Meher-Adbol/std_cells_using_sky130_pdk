**AND gate tr tf

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

Vdd vdd gnd DC 1.8
V1 a gnd pulse(0 1.8 0p 20p 20p 1n 2n) dc 0
V2 b gnd pulse(0 1.8 0p 20p 20p 2n 4n) dc 0

x1 Vdd gnd b a a Vout andg

.subckt andg vdd gnd b a a1 Vout
xm01 out b vdd vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.27 as=0.381 ad=0.381 ps=3.14 pd=3.14
xm02 out b gnd gnd sky130_fd_pr__nfet_01v8 l=0.15 w=0.42 as=0.126 ad=0.126 ps=1.44 pd=1.44

xm03 out1 out vdd vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.27 as=0.381 ad=0.381 ps=3.14 pd=3.14
xm04 out1 a vdd vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.27 as=0.381 ad=0.381 ps=3.14 pd=3.14
xm05 out1 out x gnd sky130_fd_pr__nfet_01v8 l=0.15 w=0.42 as=0.252 ad=0.252 ps=2.28 pd=2.28
xm06 x a1 gnd gnd sky130_fd_pr__nfet_01v8 l=0.15 w=0.42 as=0.252 ad=0.252 ps=2.28 pd=2.28
xm07 out1 out x gnd sky130_fd_pr__nfet_01v8 l=0.15 w=0.42 as=0.252 ad=0.252 ps=2.28 pd=2.28
xm08 x a1 gnd gnd sky130_fd_pr__nfet_01v8 l=0.15 w=0.42 as=0.252 ad=0.252 ps=2.28 pd=2.28

xm09 Vout out1 vdd vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.27 as=0.381 ad=0.381 ps=3.14 pd=3.14
xm10 Vout out1 gnd gnd sky130_fd_pr__nfet_01v8 l=0.15 w=0.42 as=0.126 ad=0.126 ps=1.44 pd=1.44
.ends

.tran 1ps 8ns 0 10p

.control 
run

meas tran tr TRIG v(Vout) VAL = 0.36 RISE = 1 TARG v(Vout) VAL = 1.44 RISE = 1 
meas tran tf TRIG v(Vout) VAL = 1.44 FALL = 2 TARG v(Vout) VAL = 0.36 FALL = 2


let delt = abs(tr - tf)
print delt
plot v(out) v(out1) v(Vout) 
.endc
